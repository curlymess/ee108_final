// This module is just a big ROM which allows you to look up the bitmap
//  for a given character.

module tcgrom(
    input [8:0] addr,
    output reg [7:0] data
);
    // A memory is implemented using a case statement 
    always @(addr)
        case (addr)
            // PLAY
            9'h000: data = 8'b00010000; // %   *         %
            9'h001: data = 8'b00011000; // %   **        %
            9'h002: data = 8'b00011100; // %   ***       %
            9'h003: data = 8'b00011110; // %   ****      %
            9'h004: data = 8'b00011110; // %   ****      %
            9'h005: data = 8'b00011100; // %   ***       %
            9'h006: data = 8'b00011000; // %   **        %
            9'h007: data = 8'b00010000; // %   *         %
            
            // PAUSE
            9'h008: data = 8'b00000000; // %             %
            9'h009: data = 8'b11100111; // %   ***  ***  %
            9'h00a: data = 8'b11100111; // %   ***  ***  %
            9'h00b: data = 8'b11100111; // %   ***  ***  %
            9'h00c: data = 8'b11100111; // %   ***  ***  %
            9'h00d: data = 8'b11100111; // %   ***  ***  %
            9'h00e: data = 8'b11100111; // %   ***  ***  %
            9'h00f: data = 8'b11100111; // %   ***  ***  %

            // NEXT
            9'h010: data = 8'b00000000; // %             %
            9'h011: data = 8'b00000100; // %       *     %
            9'h012: data = 8'b00000110; // %       **    %
            9'h013: data = 8'b01111111; // %   *******   %
            9'h014: data = 8'b01111111; // %   *******   %
            9'h015: data = 8'b00000110; // %       **    %
            9'h016: data = 8'b00000100; // %       *     %
            9'h017: data = 8'b00000000; // %             %
            
            // FAST FORWARD
            9'h018: data = 8'b00000000; // %             %
            9'h019: data = 8'b10000000; // %   *         %
            9'h01a: data = 8'b11000100; // %   **   *    %
            9'h01b: data = 8'b11100110; // %   ***  **   %
            9'h01c: data = 8'b11111111; // %   **** ***  %
            9'h01d: data = 8'b11100110; // %   ***  **   %
            9'h01e: data = 8'b11000100; // %   **   *    %
            9'h01f: data = 8'b10000000; // %   *         %
  
            // REWIND
            9'h028: data = 8'b00000000; // %             %
            9'h029: data = 8'b00000001; // %          *  %
            9'h02a: data = 8'b00100011; // %     *   **  %
            9'h02b: data = 8'b01100111; // %    **  ***  %
            9'h02c: data = 8'b11111111; // %   *** ****  %
            9'h02d: data = 8'b01100111; // %    **  ***  %
            9'h02e: data = 8'b00100011; // %     *   **  %
            9'h02f: data = 8'b00000001; // %          *  %
  
            9'h030: data = 8'b01111110; // %   ******    %
            9'h031: data = 8'b01100000; // %   **        %
            9'h032: data = 8'b01100000; // %   **        %
            9'h033: data = 8'b01111000; // %   ****      %
            9'h034: data = 8'b01100000; // %   **        %
            9'h035: data = 8'b01100000; // %   **        %
            9'h036: data = 8'b01111110; // %   ******    %
            9'h037: data = 8'b00000000; // %             %
    
            9'h038: data = 8'b00111100; // %    ****     %
            9'h039: data = 8'b01100110; // %   **  **    %
            9'h03a: data = 8'b01100000; // %   **        %
            9'h03b: data = 8'b01101110; // %   ** ***    %
            9'h03c: data = 8'b01100110; // %   **  **    %
            9'h03d: data = 8'b01100110; // %   **  **    %
            9'h03e: data = 8'b00111100; // %    ****     %
            9'h03f: data = 8'b00000000; // %             %
  
            9'h040: data = 8'b01100110; // %   **  **    %
            9'h041: data = 8'b01100110; // %   **  **    %
            9'h042: data = 8'b01100110; // %   **  **    %
            9'h043: data = 8'b01111110; // %   ******    %
            9'h044: data = 8'b01100110; // %   **  **    %
            9'h045: data = 8'b01100110; // %   **  **    %
            9'h046: data = 8'b01100110; // %   **  **    %
            9'h047: data = 8'b00000000; // %             %
  
            9'h048: data = 8'b00111100; // %    ****     %
            9'h049: data = 8'b00011000; // %     **      %
            9'h04a: data = 8'b00011000; // %     **      %
            9'h04b: data = 8'b00011000; // %     **      %
            9'h04c: data = 8'b00011000; // %     **      %
            9'h04d: data = 8'b00011000; // %     **      %
            9'h04e: data = 8'b00111100; // %    ****     %
            9'h04f: data = 8'b00000000; // %             %
  
            9'h0a0: data = 8'b01111110; // %   ******    %
            9'h0a1: data = 8'b00011000; // %     **      %
            9'h0a2: data = 8'b00011000; // %     **      %
            9'h0a3: data = 8'b00011000; // %     **      %
            9'h0a4: data = 8'b00011000; // %     **      %
            9'h0a5: data = 8'b00011000; // %     **      %
            9'h0a6: data = 8'b00011000; // %     **      %
            9'h0a7: data = 8'b00000000; // %             %
    
            9'h0b8: data = 8'b01100011; // %   **   **   %
            9'h0b9: data = 8'b01100011; // %   **   **   %
            9'h0ba: data = 8'b01100011; // %   **   **   %
            9'h0bb: data = 8'b01101011; // %   ** * **   %
            9'h0bc: data = 8'b01111111; // %   *******   %
            9'h0bd: data = 8'b01110111; // %   *** ***   %
            9'h0be: data = 8'b01100011; // %   **   **   %
            9'h0bf: data = 8'b00000000; // %             %
  
            9'h180: data = 8'b00111100; // %    ****     %
            9'h181: data = 8'b01100110; // %   **  **    %
            9'h182: data = 8'b01101110; // %   ** ***    %
            9'h183: data = 8'b01110110; // %   *** **    %
            9'h184: data = 8'b01100110; // %   **  **    %
            9'h185: data = 8'b01100110; // %   **  **    %
            9'h186: data = 8'b00111100; // %    ****     %
            9'h187: data = 8'b00000000; // %             %
  
            9'h188: data = 8'b00011000; // %     **      %
            9'h189: data = 8'b00011000; // %     **    . %
            9'h18a: data = 8'b00111000; // %    ***      %
            9'h18b: data = 8'b00011000; // %     **      %
            9'h18c: data = 8'b00011000; // %     **      %
            9'h18d: data = 8'b00011000; // %     **      %
            9'h18e: data = 8'b01111110; // %   ******    %
            9'h18f: data = 8'b00000000; // %             %
  
            9'h190: data = 8'b00111100; // %    ****     %
            9'h191: data = 8'b01100110; // %   **  **    %
            9'h192: data = 8'b00000110; // %       **    %
            9'h193: data = 8'b00001100; // %      **     %
            9'h194: data = 8'b00110000; // %    **       %
            9'h195: data = 8'b01100000; // %   **        %
            9'h196: data = 8'b01111110; // %   ******    %
            9'h197: data = 8'b00000000; // %             %
  
            9'h198: data = 8'b00111100; // %    ****     %
            9'h199: data = 8'b01100110; // %   **  **    %
            9'h19a: data = 8'b00000110; // %       **    %
            9'h19b: data = 8'b00011100; // %     ***     %
            9'h19c: data = 8'b00000110; // %       **    %
            9'h19d: data = 8'b01100110; // %   **  **    %
            9'h19e: data = 8'b00111100; // %    ****     %
            9'h19f: data = 8'b00000000; // %             %
            
            default: data = 8'd0;
        endcase

endmodule
