module sample_adder(
    input clk,
    input reset
);

endmodule